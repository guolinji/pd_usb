library verilog;
use verilog.vl_types.all;
entity tb_prl_phy_top is
end tb_prl_phy_top;
